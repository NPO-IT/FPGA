module memDblArray
(
	input reset,
	input clk,
	input iRQ,
	input [4:0]iNumRQ,
	output reg[7:0]MARK,
	output reg[7:0]m1b1,
	output reg[7:0]m1b2,
	output reg[7:0]m1b3,
	output reg[7:0]m1b4,
	output reg[7:0]m2b1,
	output reg[7:0]m2b2,
	output reg[7:0]m2b3,
	output reg[7:0]m2b4,
	output reg[7:0]m3b1,
	output reg[7:0]m3b2,
	output reg[7:0]m3b3,
	output reg[7:0]m3b4,
	output reg[7:0]CRC8,

	output reg test
);

`define WAIT 0
`define TX 1
`define DONE 2

reg [7:0] Memories [0:31][0:13] = '{
'{8'd129,	8'd130,	8'd131,	8'd132,	8'd135,	8'd136,	8'd166,	8'd50,	8'd148,	8'd149,	8'd50,	8'd50,	8'd190,	8'd186},	//rq# 0
'{8'd133,	8'd134,	8'd7,	8'd8,	8'd132,	8'd133,	8'd134,	8'd50,	8'd154,	8'd155,	8'd50,	8'd50,	8'd15,	8'd166},	//rq# 1
'{8'd9,		8'd138,	8'd139,	8'd140,	8'd129,	8'd130,	8'd131,	8'd50,	8'd129,	8'd130,	8'd50,	8'd50,	8'd170,	8'd20},		//rq# 2
'{8'd141,	8'd142,	8'd143,	8'd144,	8'd137,	8'd138,	8'd139,	8'd50,	8'd131,	8'd132,	8'd50,	8'd50,	8'd200,	8'd0},		//rq# 3
'{8'd159,	8'd160,	8'd161,	8'd162,	8'd135,	8'd136,	8'd167,	8'd50,	8'd133,	8'd134,	8'd50,	8'd50,	8'd187,	8'd198},	//rq# 4
'{8'd145,	8'd146,	8'd147,	8'd148,	8'd140,	8'd141,	8'd142,	8'd50,	8'd135,	8'd136,	8'd50,	8'd50,	8'd13,	8'd180},	//rq# 5
'{8'd149,	8'd150,	8'd151,	8'd152,	8'd143,	8'd144,	8'd145,	8'd50,	8'd137,	8'd138,	8'd50,	8'd50,	8'd79,	8'd187},	//rq# 6
'{8'd153,	8'd154,	8'd155,	8'd156,	8'd146,	8'd147,	8'd148,	8'd50,	8'd139,	8'd140,	8'd50,	8'd50,	8'd126,	8'd4},		//rq# 7
'{8'd129,	8'd130,	8'd131,	8'd132,	8'd135,	8'd136,	8'd166,	8'd50,	8'd148,	8'd149,	8'd50,	8'd50,	8'd190,	8'd186},	//rq# 8
'{8'd133,	8'd134,	8'd7,	8'd8,	8'd132,	8'd133,	8'd134,	8'd50,	8'd154,	8'd155,	8'd50,	8'd50,	8'd15,	8'd166},	//rq# 9
'{8'd9,		8'd138,	8'd139,	8'd140,	8'd149,	8'd150,	8'd151,	8'd50,	8'd141,	8'd142,	8'd50,	8'd50,	8'd72,	8'd6},		//rq# 10
'{8'd141,	8'd142,	8'd143,	8'd144,	8'd152,	8'd153,	8'd154,	8'd50,	8'd143,	8'd144,	8'd50,	8'd50,	8'd210,	8'd43},		//rq# 11
'{8'd159,	8'd160,	8'd161,	8'd162,	8'd135,	8'd136,	8'd155,	8'd50,	8'd145,	8'd146,	8'd50,	8'd50,	8'd209,	8'd92},		//rq# 12
'{8'd157,	8'd163,	8'd164,	8'd165,	8'd156,	8'd157,	8'd159,	8'd50,	8'd147,	8'd150,	8'd50,	8'd50,	8'd78,	8'd89},		//rq# 13
'{8'd166,	8'd167,	8'd168,	8'd176,	8'd160,	8'd161,	8'd162,	8'd50,	8'd151,	8'd152,	8'd50,	8'd50,	8'd119,	8'd39},		//rq# 14
'{8'd177,	8'd50,	8'd50,	8'd50,	8'd163,	8'd164,	8'd165,	8'd50,	8'd153,	8'd156,	8'd50,	8'd50,	8'd135,	8'd26},		//rq# 15
'{8'd129,	8'd130,	8'd131,	8'd132,	8'd135,	8'd136,	8'd40,	8'd50,	8'd148,	8'd149,	8'd50,	8'd50,	8'd234,	8'd57},		//rq# 16
'{8'd133,	8'd134,	8'd7,	8'd8,	8'd132,	8'd133,	8'd134,	8'd50,	8'd154,	8'd155,	8'd50,	8'd50,	8'd15,	8'd166},	//rq# 17
'{8'd9,		8'd138,	8'd139,	8'd140,	8'd176,	8'd177,	8'd50,	8'd50,	8'd31,	8'd160,	8'd50,	8'd50,	8'd195,	8'd66},		//rq# 18
'{8'd141,	8'd142,	8'd143,	8'd144,	8'd50,	8'd50,	8'd50,	8'd50,	8'd161,	8'd162,	8'd50,	8'd50,	8'd153,	8'd37},		//rq# 19
'{8'd159,	8'd160,	8'd161,	8'd162,	8'd135,	8'd136,	8'd167,	8'd50,	8'd176,	8'd177,	8'd50,	8'd50,	8'd107,	8'd95},		//rq# 20
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116},	//rq# 21
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116},	//rq# 22
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116},	//rq# 23
'{8'd129,	8'd130,	8'd131,	8'd132,	8'd135,	8'd136,	8'd166,	8'd50,	8'd148,	8'd149,	8'd50,	8'd50,	8'd190,	8'd186},	//rq# 24
'{8'd133,	8'd134,	8'd7,	8'd8,	8'd132,	8'd133,	8'd134,	8'd50,	8'd154,	8'd155,	8'd50,	8'd50,	8'd15,	8'd166},	//rq# 25
'{8'd9,		8'd138,	8'd139,	8'd140,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd1,	8'd182},	//rq# 26
'{8'd141,	8'd142,	8'd143,	8'd144,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd188,	8'd95},		//rq# 27
'{8'd159,	8'd160,	8'd161,	8'd162,	8'd135,	8'd136,	8'd178,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd96,	8'd128},	//rq# 28
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116},	//rq# 29
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116},	//rq# 30
'{8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd50,	8'd198,	8'd116}		//rq# 31
};

reg [1:0]state;


always@(posedge clk)
begin
	if (~reset) begin								// initial
		
	end else begin									// main
		case (state)
			`WAIT: begin
				if (~iRQ) state <= `TX;
			end
			`TX: begin
				MARK <= 8'b11001100;
				m1b1 <= Memories[iNumRQ][0];
				m1b2 <= Memories[iNumRQ][1];
				m1b3 <= Memories[iNumRQ][2];
				m1b4 <= Memories[iNumRQ][3];
				m2b1 <= Memories[iNumRQ][4];
				m2b2 <= Memories[iNumRQ][5];
				m2b3 <= Memories[iNumRQ][6];
				m2b4 <= Memories[iNumRQ][7];
				m3b1 <= Memories[iNumRQ][8];
				m3b2 <= Memories[iNumRQ][9];
				m3b3 <= Memories[iNumRQ][10];
				m3b4 <= Memories[iNumRQ][11];
				CRC8 <= Memories[iNumRQ][12];
			end
			`DONE: begin
				if (iRQ) state <= `WAIT;
			end
		endcase
	end
end
endmodule
